library verilog;
use verilog.vl_types.all;
entity VGA_SRAM_interface_v_unit is
end VGA_SRAM_interface_v_unit;
