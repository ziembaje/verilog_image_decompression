library verilog;
use verilog.vl_types.all;
entity UART_SRAM_interface_v_unit is
end UART_SRAM_interface_v_unit;
