library verilog;
use verilog.vl_types.all;
entity Milestone_1_v_unit is
end Milestone_1_v_unit;
