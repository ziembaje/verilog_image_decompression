library verilog;
use verilog.vl_types.all;
entity UART_Receive_Controller_v_unit is
end UART_Receive_Controller_v_unit;
