library verilog;
use verilog.vl_types.all;
entity final_project_v_unit is
end final_project_v_unit;
